library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.ALL;

entity Distribute is
    port (
		  CLK : in  STD_LOGIC;
		  
		  byte_in : in  STD_LOGIC := '0';
		  q_in : in STD_LOGIC_VECTOR (7 downto 0);
		  swap_out : out  STD_LOGIC := '0';
		  set_out : out STD_LOGIC := '0';
		  multiplex_out : out STD_LOGIC := '0';
		  data_out: out STD_LOGIC_VECTOR (7 downto 0); 
		  address : out std_logic_vector(8 downto 0); --400 addresses
		  
		  debug_swap : out STD_LOGIC := '0';
		  debug_reset : out STD_LOGIC := '0';
		  debug_onShiftClocks : out STD_LOGIC := '1'
	 );
end Distribute;

architecture Behavioral of Distribute is

type T_PHASE_CORRECTION is array (0 to 399) of integer range 0 to 255;
	constant PHASE_CORRECTION : T_PHASE_CORRECTION := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
																		0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
		
	 signal s_boardEnable : STD_LOGIC := '1';
	 signal s_ByteCounter : integer range 0 to 399 := 0;
	  
	 signal s_data_out : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	 signal s_address : std_logic_vector(8 downto 0) := (others => '0');
	 signal s_swap_out :  STD_LOGIC := '0';
	 signal s_set_out : STD_LOGIC := '0';
	 
	 signal s_debug_swap : STD_LOGIC := '0';
	 signal s_debug_onShiftClocks : STD_LOGIC := '1';
begin
    Distribute: process (clk) begin
        if (rising_edge(clk)) then
				if (byte_in = '1') then --a byte of data is ready
					
					if (q_in = "11111110" AND s_boardEnable = '1') then --254 is start phases
						s_ByteCounter <= 0;
						s_swap_out <= '0';
						s_set_out <= '0';
					elsif (q_in = "11111101") then --253 is swap
						s_debug_swap <= not s_debug_swap;
						s_set_out <= '0';
						s_swap_out <= '1';
						s_ByteCounter <= 0;
						
					elsif (q_in = "10010110") then --150 is switch off clocks
						s_debug_onShiftClocks <= '0';
					elsif (q_in = "10010111") then --151 is switch on clocks
						s_debug_onShiftClocks <= '1';
						
					elsif (q_in = "11000000") then --192 board primary
						s_boardEnable <= '1';
					elsif (q_in = "11000001") then --193 board secondary
						s_boardEnable <= '0';
						
					elsif (s_boardEnable = '1') then-- any other byte is for the delay lines. send only if the board is enabled
						--s_data_out <= q_in;
						s_address <= std_logic_vector(to_unsigned(s_ByteCounter, 9));
						s_swap_out <= '0';
						s_set_out <= '1';
						s_ByteCounter <= s_ByteCounter + 1;
						
						if (q_in = "00100000") then
							s_data_out <= q_in; -- a phase of 32 represents "off" so no phase correction
						else
							s_data_out <= std_logic_vector( to_unsigned( to_integer(unsigned(q_in)) + PHASE_CORRECTION(s_ByteCounter), 8 ) ) and "00011111";
						end if;
						
					end if;
				else
					s_swap_out <= '0';
					s_set_out <= '0';
				end if;
				
				
		  end if;
 end process;
 debug_swap <= s_debug_swap;
 debug_reset <= s_boardEnable;
 debug_onShiftClocks <= s_debug_onShiftClocks;
 
 data_out <= s_data_out;
 address <= s_address;
 swap_out <= s_swap_out;
 set_out <= s_set_out;
 
end Behavioral;
